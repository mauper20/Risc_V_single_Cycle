
/******************************************************************
* Description
*	and logica
*	1.0
* Author:
*	Adrian Guevara, Mauricio Peralta
* email:
*	mperalta.osorio@iteso.mx
* Date:
*	25/10/2021
******************************************************************/
module ORGate
(
	input A,
	input B,
	output C
);


assign C = A | B;

endmodule